library verilog;
use verilog.vl_types.all;
entity my_package_vlg_vec_tst is
end my_package_vlg_vec_tst;
